module top_module( output one );

// Insert your code here
    wire x;
    assign one = 1'b1;
    ddasa

endmodule